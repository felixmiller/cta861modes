
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package video_timings_pkg is

    type video_timing_r is record
        name        : string(1 to 20);
        vic         : natural range 0 to 255;
        pxl_clk_khz : natural range 0 to 2**13-1;
        interlaced  : boolean;
        dbl_clkd    : boolean;
        hactive     : natural range 0 to 2**13-1;
        vactive     : natural range 0 to 2**13-1;
        hfront      : natural range 0 to 2**13-1;
        hsync       : natural range 0 to 2**13-1;
        hback       : natural range 0 to 2**13-1;
        hpol        : std_logic;
        vfront      : natural range 0 to 2**13-1;
        vsync       : natural range 0 to 2**13-1;
        vback       : natural range 0 to 2**13-1;
        vpol        : std_logic;
        ln          : integer range 0 to 7;
    end record;

    type video_timings_a is array (0 to 219) of video_timing_r;

    constant video_timings : video_timings_a := (
    --  VIC    |  Name              | VIC | Pixel Clk kHz | interlaced | double clocked | hactive | vactive | hfront | hsync | hback | hpol | vfront | vsync | vback | vpol | ln

          1 => ("640x480@60Hz        ",    1,          25175,       false,           false,      640,      480,      16,     96,     48,   '0',      10,      2,     33,   '0',  1 ),
          2 => ("720x480@60Hz        ",    2,          27000,       false,           false,      720,      480,      16,     62,     60,   '0',       9,      6,     30,   '0',  7 ),
          3 => ("720x480@60Hz        ",    3,          27000,       false,           false,      720,      480,      16,     62,     60,   '0',       9,      6,     30,   '0',  7 ),
          4 => ("1280x720@60Hz       ",    4,          74250,       false,           false,     1280,      720,     110,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
          5 => ("1920x1080i@60Hz     ",    5,          74250,        true,           false,     1920,     1080,      88,     44,    148,   '1',       4,     10,     31,   '1',  1 ),
          6 => ("720x480i@60Hz       ",    6,          13500,        true,            true,      720,      480,      19,     62,     57,   '0',       8,      6,     31,   '0',  4 ),
          7 => ("720x480i@60Hz       ",    7,          13500,        true,            true,      720,      480,      19,     62,     57,   '0',       8,      6,     31,   '0',  4 ),
          8 => ("720x240@60Hz        ",    8,          13500,       false,            true,      720,      240,      19,     62,     57,   '0',       4,      3,     15,   '0',  4 ),
          9 => ("720x240@60Hz        ",    9,          13500,       false,            true,      720,      240,      19,     62,     57,   '0',       4,      3,     15,   '0',  4 ),
         10 => ("2880x480i@60Hz      ",   10,          54000,        true,           false,     2880,      480,      76,    248,    228,   '0',       8,      6,     31,   '0',  4 ),
         11 => ("2880x480i@60Hz      ",   11,          54000,        true,           false,     2880,      480,      76,    248,    228,   '0',       8,      6,     31,   '0',  4 ),
         12 => ("2880x240@60Hz       ",   12,          54000,       false,           false,     2880,      240,      76,    248,    228,   '0',       4,      3,     15,   '0',  4 ),
         13 => ("2880x240@60Hz       ",   13,          54000,       false,           false,     2880,      240,      76,    248,    228,   '0',       4,      3,     15,   '0',  4 ),
         14 => ("1440x480@60Hz       ",   14,          54000,       false,           false,     1440,      480,      32,    124,    120,   '0',       9,      6,     30,   '0',  7 ),
         15 => ("1440x480@60Hz       ",   15,          54000,       false,           false,     1440,      480,      32,    124,    120,   '0',       9,      6,     30,   '0',  7 ),
         16 => ("1920x1080@60Hz      ",   16,         148500,       false,           false,     1920,     1080,      88,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         17 => ("720x576@50Hz        ",   17,          27000,       false,           false,      720,      576,      12,     64,     68,   '0',       5,      5,     39,   '0',  1 ),
         18 => ("720x576@50Hz        ",   18,          27000,       false,           false,      720,      576,      12,     64,     68,   '0',       5,      5,     39,   '0',  1 ),
         19 => ("1280x720@50Hz       ",   19,          74250,       false,           false,     1280,      720,     440,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         20 => ("1920x1080i@50Hz     ",   20,          74250,        true,           false,     1920,     1080,     528,     44,    148,   '1',       4,     10,     31,   '1',  1 ),
         21 => ("720x576i@50Hz       ",   21,          13500,        true,            true,      720,      576,      12,     63,     69,   '0',       4,      6,     39,   '0',  1 ),
         22 => ("720x576i@50Hz       ",   22,          13500,        true,            true,      720,      576,      12,     63,     69,   '0',       4,      6,     39,   '0',  1 ),
         23 => ("720x288@50Hz        ",   23,          13500,       false,            true,      720,      288,      12,     63,     69,   '0',       2,      3,     19,   '0',  1 ),
         24 => ("720x288@50Hz        ",   24,          13500,       false,            true,      720,      288,      12,     63,     69,   '0',       2,      3,     19,   '0',  1 ),
         25 => ("2880x576i@50Hz      ",   25,          54000,        true,           false,     2880,      576,      48,    252,    276,   '0',       4,      6,     39,   '0',  1 ),
         26 => ("2880x576i@50Hz      ",   26,          54000,        true,           false,     2880,      576,      48,    252,    276,   '0',       4,      6,     39,   '0',  1 ),
         27 => ("2880x288@50Hz       ",   27,          54000,       false,           false,     2880,      288,      48,    252,    276,   '0',       2,      3,     19,   '0',  1 ),
         28 => ("2880x288@50Hz       ",   28,          54000,       false,           false,     2880,      288,      48,    252,    276,   '0',       2,      3,     19,   '0',  1 ),
         29 => ("1440x576@50Hz       ",   29,          54000,       false,           false,     1440,      576,      24,    128,    136,   '0',       5,      5,     39,   '0',  1 ),
         30 => ("1440x576@50Hz       ",   30,          54000,       false,           false,     1440,      576,      24,    128,    136,   '0',       5,      5,     39,   '0',  1 ),
         31 => ("1920x1080@50Hz      ",   31,         148500,       false,           false,     1920,     1080,     528,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         32 => ("1920x1080@24Hz      ",   32,          74250,       false,           false,     1920,     1080,     638,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         33 => ("1920x1080@25Hz      ",   33,          74250,       false,           false,     1920,     1080,     528,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         34 => ("1920x1080@30Hz      ",   34,          74250,       false,           false,     1920,     1080,      88,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         35 => ("2880x480@60Hz       ",   35,         108000,       false,           false,     2880,      480,      64,    248,    240,   '0',       9,      6,     30,   '0',  7 ),
         36 => ("2880x480@60Hz       ",   36,         108000,       false,           false,     2880,      480,      64,    248,    240,   '0',       9,      6,     30,   '0',  7 ),
         37 => ("2880x576@50Hz       ",   37,         108000,       false,           false,     2880,      576,      48,    256,    272,   '0',       5,      5,     39,   '0',  1 ),
         38 => ("2880x576@50Hz       ",   38,         108000,       false,           false,     2880,      576,      48,    256,    272,   '0',       5,      5,     39,   '0',  1 ),
         39 => ("1920x1080i@50Hz     ",   39,          72000,        true,           false,     1920,     1080,      32,    168,    184,   '1',      46,     10,    114,   '0',  1 ),
         40 => ("1920x1080i@100Hz    ",   40,         148500,        true,           false,     1920,     1080,     528,     44,    148,   '1',       4,     10,     31,   '1',  1 ),
         41 => ("1280x720@100Hz      ",   41,         148500,       false,           false,     1280,      720,     440,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         42 => ("720x576@100Hz       ",   42,          54000,       false,           false,      720,      576,      12,     64,     68,   '0',       5,      5,     39,   '0',  1 ),
         43 => ("720x576@100Hz       ",   43,          54000,       false,           false,      720,      576,      12,     64,     68,   '0',       5,      5,     39,   '0',  1 ),
         44 => ("720x576i@100Hz      ",   44,          27000,        true,            true,      720,      576,      12,     63,     69,   '0',       4,      6,     39,   '0',  1 ),
         45 => ("720x576i@100Hz      ",   45,          27000,        true,            true,      720,      576,      12,     63,     69,   '0',       4,      6,     39,   '0',  1 ),
         46 => ("1920x1080i@120Hz    ",   46,         148500,        true,           false,     1920,     1080,      88,     44,    148,   '1',       4,     10,     31,   '1',  1 ),
         47 => ("1280x720@120Hz      ",   47,         148500,       false,           false,     1280,      720,     110,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         48 => ("720x480@120Hz       ",   48,          54000,       false,           false,      720,      480,      16,     62,     60,   '0',       9,      6,     30,   '0',  7 ),
         49 => ("720x480@120Hz       ",   49,          54000,       false,           false,      720,      480,      16,     62,     60,   '0',       9,      6,     30,   '0',  7 ),
         50 => ("720x480i@120Hz      ",   50,          27000,        true,            true,      720,      480,      19,     62,     57,   '0',       8,      6,     31,   '0',  4 ),
         51 => ("720x480i@120Hz      ",   51,          27000,        true,            true,      720,      480,      19,     62,     57,   '0',       8,      6,     31,   '0',  4 ),
         52 => ("720x576@200Hz       ",   52,         108000,       false,           false,      720,      576,      12,     64,     68,   '0',       5,      5,     39,   '0',  1 ),
         53 => ("720x576@200Hz       ",   53,         108000,       false,           false,      720,      576,      12,     64,     68,   '0',       5,      5,     39,   '0',  1 ),
         54 => ("720x576i@200Hz      ",   54,          54000,        true,            true,      720,      576,      12,     63,     69,   '0',       4,      6,     39,   '0',  1 ),
         55 => ("720x576i@200Hz      ",   55,          54000,        true,            true,      720,      576,      12,     63,     69,   '0',       4,      6,     39,   '0',  1 ),
         56 => ("720x480@240Hz       ",   56,         108000,       false,           false,      720,      480,      16,     62,     60,   '0',       9,      6,     30,   '0',  7 ),
         57 => ("720x480@240Hz       ",   57,         108000,       false,           false,      720,      480,      16,     62,     60,   '0',       9,      6,     30,   '0',  7 ),
         58 => ("720x480i@240Hz      ",   58,          54000,        true,            true,      720,      480,      19,     62,     57,   '0',       8,      6,     31,   '0',  4 ),
         59 => ("720x480i@240Hz      ",   59,          54000,        true,            true,      720,      480,      19,     62,     57,   '0',       8,      6,     31,   '0',  4 ),
         60 => ("1280x720@24Hz       ",   60,          59400,       false,           false,     1280,      720,    1760,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         61 => ("1280x720@25Hz       ",   61,          74250,       false,           false,     1280,      720,    2420,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         62 => ("1280x720@30Hz       ",   62,          74250,       false,           false,     1280,      720,    1760,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         63 => ("1920x1080@120Hz     ",   63,         297000,       false,           false,     1920,     1080,      88,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         64 => ("1920x1080@100Hz     ",   64,         297000,       false,           false,     1920,     1080,     528,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         65 => ("1280x720@24Hz       ",   65,          59400,       false,           false,     1280,      720,    1760,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         66 => ("1280x720@25Hz       ",   66,          74250,       false,           false,     1280,      720,    2420,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         67 => ("1280x720@30Hz       ",   67,          74250,       false,           false,     1280,      720,    1760,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         68 => ("1280x720@50Hz       ",   68,          74250,       false,           false,     1280,      720,     440,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         69 => ("1280x720@60Hz       ",   69,          74250,       false,           false,     1280,      720,     110,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         70 => ("1280x720@100Hz      ",   70,         148500,       false,           false,     1280,      720,     440,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         71 => ("1280x720@120Hz      ",   71,         148500,       false,           false,     1280,      720,     110,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         72 => ("1920x1080@24Hz      ",   72,          74250,       false,           false,     1920,     1080,     638,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         73 => ("1920x1080@25Hz      ",   73,          74250,       false,           false,     1920,     1080,     528,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         74 => ("1920x1080@30Hz      ",   74,          74250,       false,           false,     1920,     1080,      88,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         75 => ("1920x1080@50Hz      ",   75,         148500,       false,           false,     1920,     1080,     528,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         76 => ("1920x1080@60Hz      ",   76,         148500,       false,           false,     1920,     1080,      88,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         77 => ("1920x1080@100Hz     ",   77,         297000,       false,           false,     1920,     1080,     528,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         78 => ("1920x1080@120Hz     ",   78,         297000,       false,           false,     1920,     1080,      88,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         79 => ("1680x720@24Hz       ",   79,          59400,       false,           false,     1680,      720,    1360,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         80 => ("1680x720@25Hz       ",   80,          59400,       false,           false,     1680,      720,    1228,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         81 => ("1680x720@30Hz       ",   81,          59400,       false,           false,     1680,      720,     700,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         82 => ("1680x720@50Hz       ",   82,          82500,       false,           false,     1680,      720,     260,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         83 => ("1680x720@60Hz       ",   83,          99000,       false,           false,     1680,      720,     260,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
         84 => ("1680x720@100Hz      ",   84,         165000,       false,           false,     1680,      720,      60,     40,    220,   '1',       5,      5,     95,   '1',  1 ),
         85 => ("1680x720@120Hz      ",   85,         198000,       false,           false,     1680,      720,      60,     40,    220,   '1',       5,      5,     95,   '1',  1 ),
         86 => ("2560x1080@24Hz      ",   86,          99000,       false,           false,     2560,     1080,     998,     44,    148,   '1',       4,      5,     11,   '1',  1 ),
         87 => ("2560x1080@25Hz      ",   87,          90000,       false,           false,     2560,     1080,     448,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         88 => ("2560x1080@30Hz      ",   88,         118800,       false,           false,     2560,     1080,     768,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         89 => ("2560x1080@50Hz      ",   89,         185625,       false,           false,     2560,     1080,     548,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
         90 => ("2560x1080@60Hz      ",   90,         198000,       false,           false,     2560,     1080,     248,     44,    148,   '1',       4,      5,     11,   '1',  1 ),
         91 => ("2560x1080@100Hz     ",   91,         371250,       false,           false,     2560,     1080,     218,     44,    148,   '1',       4,      5,    161,   '1',  1 ),
         92 => ("2560x1080@120Hz     ",   92,         495000,       false,           false,     2560,     1080,     548,     44,    148,   '1',       4,      5,    161,   '1',  1 ),
         93 => ("3840x2160@24Hz      ",   93,         297000,       false,           false,     3840,     2160,    1276,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
         94 => ("3840x2160@25Hz      ",   94,         297000,       false,           false,     3840,     2160,    1056,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
         95 => ("3840x2160@30Hz      ",   95,         297000,       false,           false,     3840,     2160,     176,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
         96 => ("3840x2160@50Hz      ",   96,         594000,       false,           false,     3840,     2160,    1056,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
         97 => ("3840x2160@60Hz      ",   97,         594000,       false,           false,     3840,     2160,     176,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
         98 => ("4096x2160@24Hz      ",   98,         297000,       false,           false,     4096,     2160,    1020,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
         99 => ("4096x2160@25Hz      ",   99,         297000,       false,           false,     4096,     2160,     968,     88,    128,   '1',       8,     10,     72,   '1',  1 ),
        100 => ("4096x2160@30Hz      ",  100,         297000,       false,           false,     4096,     2160,      88,     88,    128,   '1',       8,     10,     72,   '1',  1 ),
        101 => ("4096x2160@50Hz      ",  101,         594000,       false,           false,     4096,     2160,     968,     88,    128,   '1',       8,     10,     72,   '1',  1 ),
        102 => ("4096x2160@60Hz      ",  102,         594000,       false,           false,     4096,     2160,      88,     88,    128,   '1',       8,     10,     72,   '1',  1 ),
        103 => ("3840x2160@24Hz      ",  103,         297000,       false,           false,     3840,     2160,    1276,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        104 => ("3840x2160@25Hz      ",  104,         297000,       false,           false,     3840,     2160,    1056,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        105 => ("3840x2160@30Hz      ",  105,         297000,       false,           false,     3840,     2160,     176,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        106 => ("3840x2160@50Hz      ",  106,         594000,       false,           false,     3840,     2160,    1056,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        107 => ("3840x2160@60Hz      ",  107,         594000,       false,           false,     3840,     2160,     176,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        108 => ("1280x720@48Hz       ",  108,          90000,       false,           false,     1280,      720,     960,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
        109 => ("1280x720@48Hz       ",  109,          90000,       false,           false,     1280,      720,     960,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
        110 => ("1680x720@48Hz       ",  110,          99000,       false,           false,     1680,      720,     810,     40,    220,   '1',       5,      5,     20,   '1',  1 ),
        111 => ("1920x1080@48Hz      ",  111,         148500,       false,           false,     1920,     1080,     638,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
        112 => ("1920x1080@48Hz      ",  112,         148500,       false,           false,     1920,     1080,     638,     44,    148,   '1',       4,      5,     36,   '1',  1 ),
        113 => ("2560x1080@48Hz      ",  113,         198000,       false,           false,     2560,     1080,     998,     44,    148,   '1',       4,      5,     11,   '1',  1 ),
        114 => ("3840x2160@48Hz      ",  114,         594000,       false,           false,     3840,     2160,    1276,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        115 => ("4096x2160@48Hz      ",  115,         594000,       false,           false,     4096,     2160,    1020,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        116 => ("3840x2160@48Hz      ",  116,         594000,       false,           false,     3840,     2160,    1276,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        117 => ("3840x2160@100Hz     ",  117,        1188000,       false,           false,     3840,     2160,    1056,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        118 => ("3840x2160@120Hz     ",  118,        1188000,       false,           false,     3840,     2160,     176,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        119 => ("3840x2160@100Hz     ",  119,        1188000,       false,           false,     3840,     2160,    1056,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        120 => ("3840x2160@120Hz     ",  120,        1188000,       false,           false,     3840,     2160,     176,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        121 => ("5120x2160@24Hz      ",  121,         396000,       false,           false,     5120,     2160,    1996,     88,    296,   '1',       8,     10,     22,   '1',  1 ),
        122 => ("5120x2160@25Hz      ",  122,         396000,       false,           false,     5120,     2160,    1696,     88,    296,   '1',       8,     10,     22,   '1',  1 ),
        123 => ("5120x2160@30Hz      ",  123,         396000,       false,           false,     5120,     2160,     664,     88,    128,   '1',       8,     10,     22,   '1',  1 ),
        124 => ("5120x2160@48Hz      ",  124,         742500,       false,           false,     5120,     2160,     746,     88,    296,   '1',       8,     10,    297,   '1',  1 ),
        125 => ("5120x2160@50Hz      ",  125,         742500,       false,           false,     5120,     2160,    1096,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        126 => ("5120x2160@60Hz      ",  126,         742500,       false,           false,     5120,     2160,     164,     88,    128,   '1',       8,     10,     72,   '1',  1 ),
        127 => ("5120x2160@100Hz     ",  127,        1485000,       false,           false,     5120,     2160,    1096,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        193 => ("5120x2160@120Hz     ",  193,        1485000,       false,           false,     5120,     2160,     164,     88,    128,   '1',       8,     10,     72,   '1',  1 ),
        194 => ("7680x4320@24Hz      ",  194,        1188000,       false,           false,     7680,     4320,    2552,    176,    592,   '1',      16,     20,    144,   '1',  1 ),
        195 => ("7680x4320@25Hz      ",  195,        1188000,       false,           false,     7680,     4320,    2352,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        196 => ("7680x4320@30Hz      ",  196,        1188000,       false,           false,     7680,     4320,     552,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        197 => ("7680x4320@48Hz      ",  197,        2376000,       false,           false,     7680,     4320,    2552,    176,    592,   '1',      16,     20,    144,   '1',  1 ),
        198 => ("7680x4320@50Hz      ",  198,        2376000,       false,           false,     7680,     4320,    2352,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        199 => ("7680x4320@60Hz      ",  199,        2376000,       false,           false,     7680,     4320,     552,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        200 => ("7680x4320@100Hz     ",  200,        4752000,       false,           false,     7680,     4320,    2112,    176,    592,   '1',      16,     20,    144,   '1',  1 ),
        201 => ("7680x4320@120Hz     ",  201,        4752000,       false,           false,     7680,     4320,     352,    176,    592,   '1',      16,     20,    144,   '1',  1 ),
        202 => ("7680x4320@24Hz      ",  202,        1188000,       false,           false,     7680,     4320,    2552,    176,    592,   '1',      16,     20,    144,   '1',  1 ),
        203 => ("7680x4320@25Hz      ",  203,        1188000,       false,           false,     7680,     4320,    2352,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        204 => ("7680x4320@30Hz      ",  204,        1188000,       false,           false,     7680,     4320,     552,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        205 => ("7680x4320@48Hz      ",  205,        2376000,       false,           false,     7680,     4320,    2552,    176,    592,   '1',      16,     20,    144,   '1',  1 ),
        206 => ("7680x4320@50Hz      ",  206,        2376000,       false,           false,     7680,     4320,    2352,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        207 => ("7680x4320@60Hz      ",  207,        2376000,       false,           false,     7680,     4320,     552,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        208 => ("7680x4320@100Hz     ",  208,        4752000,       false,           false,     7680,     4320,    2112,    176,    592,   '1',      16,     20,    144,   '1',  1 ),
        209 => ("7680x4320@120Hz     ",  209,        4752000,       false,           false,     7680,     4320,     352,    176,    592,   '1',      16,     20,    144,   '1',  1 ),
        210 => ("10240x4320@24Hz     ",  210,        1485000,       false,           false,    10240,     4320,    1492,    176,    592,   '1',      16,     20,    594,   '1',  1 ),
        211 => ("10240x4320@25Hz     ",  211,        1485000,       false,           false,    10240,     4320,    2492,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        212 => ("10240x4320@30Hz     ",  212,        1485000,       false,           false,    10240,     4320,     288,    176,    296,   '1',      16,     20,    144,   '1',  1 ),
        213 => ("10240x4320@48Hz     ",  213,        2970000,       false,           false,    10240,     4320,    1492,    176,    592,   '1',      16,     20,    594,   '1',  1 ),
        214 => ("10240x4320@50Hz     ",  214,        2970000,       false,           false,    10240,     4320,    2492,    176,    592,   '1',      16,     20,     44,   '1',  1 ),
        215 => ("10240x4320@60Hz     ",  215,        2970000,       false,           false,    10240,     4320,     288,    176,    296,   '1',      16,     20,    144,   '1',  1 ),
        216 => ("10240x4320@100Hz    ",  216,        5940000,       false,           false,    10240,     4320,    2192,    176,    592,   '1',      16,     20,    144,   '1',  1 ),
        217 => ("10240x4320@120Hz    ",  217,        5940000,       false,           false,    10240,     4320,     288,    176,    296,   '1',      16,     20,    144,   '1',  1 ),
        218 => ("4096x2160@100Hz     ",  218,        1188000,       false,           false,     4096,     2160,     800,     88,    296,   '1',       8,     10,     72,   '1',  1 ),
        219 => ("4096x2160@120Hz     ",  219,        1188000,       false,           false,     4096,     2160,      88,     88,    128,   '1',       8,     10,     72,   '1',  1 ),
     others => ("--------------------",    0,              0,       false,           false,        0,        0,       0,      0,      0,   '0',       0,      0,      0,   '0',  0 )
    );
end package video_timings_pkg;
